-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Tue Nov 29 23:18:47 2022

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY maquina_de_estados IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        X : IN STD_LOGIC := '0';
        z4 : OUT STD_LOGIC;
        z3 : OUT STD_LOGIC;
        z2 : OUT STD_LOGIC;
        z1 : OUT STD_LOGIC
    );
END maquina_de_estados;

ARCHITECTURE BEHAVIOR OF maquina_de_estados IS
    TYPE type_fstate IS (A,B,C,D,E,F,G);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,X)
    BEGIN
        IF (reset='0') THEN
            reg_fstate <= A;
            z4 <= '0';
            z3 <= '0';
            z2 <= '0';
            z1 <= '0';
        ELSE
            z4 <= '0';
            z3 <= '0';
            z2 <= '0';
            z1 <= '0';
            CASE fstate IS
                WHEN A =>
                    IF ((X = '0')) THEN
                        reg_fstate <= B;
                    ELSIF ((X = '1')) THEN
                        reg_fstate <= E;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= A;
                    END IF;

                    z4 <= '0';

                    z3 <= '0';

                    z2 <= '0';

                    z1 <= '0';
                WHEN B =>
                    reg_fstate <= C;

                    z4 <= '0';

                    z3 <= '1';

                    z2 <= '1';

                    z1 <= '0';
                WHEN C =>
                    IF ((X = '0')) THEN
                        reg_fstate <= D;
                    ELSIF ((X = '1')) THEN
                        reg_fstate <= G;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= C;
                    END IF;

                    z4 <= '1';

                    z3 <= '1';

                    z2 <= '1';

                    z1 <= '1';
                WHEN D =>
                    reg_fstate <= A;

                    z4 <= '1';

                    z3 <= '0';

                    z2 <= '0';

                    z1 <= '1';
                WHEN E =>
                    reg_fstate <= F;

                    z4 <= '1';

                    z3 <= '0';

                    z2 <= '0';

                    z1 <= '0';
                WHEN F =>
                    reg_fstate <= C;

                    z4 <= '1';

                    z3 <= '1';

                    z2 <= '0';

                    z1 <= '0';
                WHEN G =>
                    reg_fstate <= A;

                    z4 <= '1';

                    z3 <= '1';

                    z2 <= '0';

                    z1 <= '0';
                WHEN OTHERS => 
                    z4 <= 'X';
                    z3 <= 'X';
                    z2 <= 'X';
                    z1 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
